module AND(
	data1_i,
	data2_i,
	and_o
);

input data1_i, data2_i;
output and_o;

assign and_o = data1_i & data2_i;

endmodule