module IF_ID
(
    clk_i,
	flush_i,
	hazard_i,
    pc_i,
	inst_i,
    pc_o,
	inst_o
);
